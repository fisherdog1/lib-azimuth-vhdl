entity
--pasteme entity_name\
is
	port (
		);
end entity;

architecture rtl of
--pasteme entity_name\
is

begin

end architecture;
