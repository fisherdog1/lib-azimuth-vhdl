package
--pasteme package_name\
is

end package;

package body
--pasteme package_name\
is

end package body;
